module sigmoid_lut #(
    parameter WIDTH = 12,
    parameter FRAC_BITS = 6,
    parameter LUT_SIZE = 384, // Size of the LUT
    parameter ADDR_WIDTH = 9   // Address width for the LUT (log2(LUT_SIZE))
) (
    input [ADDR_WIDTH-1:0] in,
    output [WIDTH-1:0] out
);

// Sigmoid LUT values for range [0,6] in S1.5.6 format (sign-magnitude)
reg [WIDTH-1:0] lut [0:LUT_SIZE-1];

initial begin
    lut[0] = 12'd32; // x=0.0000, y=0.500000
    lut[1] = 12'd32; // x=0.0157, y=0.503916
    lut[2] = 12'd33; // x=0.0313, y=0.507832
    lut[3] = 12'd33; // x=0.0470, y=0.511747
    lut[4] = 12'd33; // x=0.0627, y=0.515661
    lut[5] = 12'd33; // x=0.0783, y=0.519572
    lut[6] = 12'd34; // x=0.0940, y=0.523481
    lut[7] = 12'd34; // x=0.1097, y=0.527388
    lut[8] = 12'd34; // x=0.1253, y=0.531291
    lut[9] = 12'd34; // x=0.1410, y=0.535190
    lut[10] = 12'd35; // x=0.1567, y=0.539085
    lut[11] = 12'd35; // x=0.1723, y=0.542975
    lut[12] = 12'd35; // x=0.1880, y=0.546859
    lut[13] = 12'd35; // x=0.2037, y=0.550739
    lut[14] = 12'd35; // x=0.2193, y=0.554612
    lut[15] = 12'd36; // x=0.2350, y=0.558478
    lut[16] = 12'd36; // x=0.2507, y=0.562337
    lut[17] = 12'd36; // x=0.2663, y=0.566189
    lut[18] = 12'd36; // x=0.2820, y=0.570033
    lut[19] = 12'd37; // x=0.2977, y=0.573868
    lut[20] = 12'd37; // x=0.3133, y=0.577694
    lut[21] = 12'd37; // x=0.3290, y=0.581512
    lut[22] = 12'd37; // x=0.3446, y=0.585319
    lut[23] = 12'd38; // x=0.3603, y=0.589116
    lut[24] = 12'd38; // x=0.3760, y=0.592903
    lut[25] = 12'd38; // x=0.3916, y=0.596679
    lut[26] = 12'd38; // x=0.4073, y=0.600443
    lut[27] = 12'd39; // x=0.4230, y=0.604195
    lut[28] = 12'd39; // x=0.4386, y=0.607935
    lut[29] = 12'd39; // x=0.4543, y=0.611663
    lut[30] = 12'd39; // x=0.4700, y=0.615378
    lut[31] = 12'd40; // x=0.4856, y=0.619079
    lut[32] = 12'd40; // x=0.5013, y=0.622766
    lut[33] = 12'd40; // x=0.5170, y=0.626439
    lut[34] = 12'd40; // x=0.5326, y=0.630098
    lut[35] = 12'd41; // x=0.5483, y=0.633742
    lut[36] = 12'd41; // x=0.5640, y=0.637370
    lut[37] = 12'd41; // x=0.5796, y=0.640983
    lut[38] = 12'd41; // x=0.5953, y=0.644580
    lut[39] = 12'd41; // x=0.6110, y=0.648161
    lut[40] = 12'd42; // x=0.6266, y=0.651725
    lut[41] = 12'd42; // x=0.6423, y=0.655273
    lut[42] = 12'd42; // x=0.6580, y=0.658803
    lut[43] = 12'd42; // x=0.6736, y=0.662315
    lut[44] = 12'd43; // x=0.6893, y=0.665810
    lut[45] = 12'd43; // x=0.7050, y=0.669287
    lut[46] = 12'd43; // x=0.7206, y=0.672745
    lut[47] = 12'd43; // x=0.7363, y=0.676185
    lut[48] = 12'd43; // x=0.7520, y=0.679605
    lut[49] = 12'd44; // x=0.7676, y=0.683007
    lut[50] = 12'd44; // x=0.7833, y=0.686389
    lut[51] = 12'd44; // x=0.7990, y=0.689751
    lut[52] = 12'd44; // x=0.8146, y=0.693093
    lut[53] = 12'd45; // x=0.8303, y=0.696416
    lut[54] = 12'd45; // x=0.8460, y=0.699718
    lut[55] = 12'd45; // x=0.8616, y=0.702999
    lut[56] = 12'd45; // x=0.8773, y=0.706259
    lut[57] = 12'd45; // x=0.8930, y=0.709499
    lut[58] = 12'd46; // x=0.9086, y=0.712717
    lut[59] = 12'd46; // x=0.9243, y=0.715914
    lut[60] = 12'd46; // x=0.9399, y=0.719089
    lut[61] = 12'd46; // x=0.9556, y=0.722243
    lut[62] = 12'd46; // x=0.9713, y=0.725374
    lut[63] = 12'd47; // x=0.9869, y=0.728484
    lut[64] = 12'd47; // x=1.0026, y=0.731572
    lut[65] = 12'd47; // x=1.0183, y=0.734637
    lut[66] = 12'd47; // x=1.0339, y=0.737680
    lut[67] = 12'd47; // x=1.0496, y=0.740700
    lut[68] = 12'd48; // x=1.0653, y=0.743697
    lut[69] = 12'd48; // x=1.0809, y=0.746672
    lut[70] = 12'd48; // x=1.0966, y=0.749624
    lut[71] = 12'd48; // x=1.1123, y=0.752552
    lut[72] = 12'd48; // x=1.1279, y=0.755458
    lut[73] = 12'd49; // x=1.1436, y=0.758341
    lut[74] = 12'd49; // x=1.1593, y=0.761200
    lut[75] = 12'd49; // x=1.1749, y=0.764036
    lut[76] = 12'd49; // x=1.1906, y=0.766848
    lut[77] = 12'd49; // x=1.2063, y=0.769638
    lut[78] = 12'd49; // x=1.2219, y=0.772403
    lut[79] = 12'd50; // x=1.2376, y=0.775146
    lut[80] = 12'd50; // x=1.2533, y=0.777864
    lut[81] = 12'd50; // x=1.2689, y=0.780559
    lut[82] = 12'd50; // x=1.2846, y=0.783231
    lut[83] = 12'd50; // x=1.3003, y=0.785879
    lut[84] = 12'd50; // x=1.3159, y=0.788503
    lut[85] = 12'd51; // x=1.3316, y=0.791104
    lut[86] = 12'd51; // x=1.3473, y=0.793681
    lut[87] = 12'd51; // x=1.3629, y=0.796235
    lut[88] = 12'd51; // x=1.3786, y=0.798764
    lut[89] = 12'd51; // x=1.3943, y=0.801271
    lut[90] = 12'd51; // x=1.4099, y=0.803754
    lut[91] = 12'd52; // x=1.4256, y=0.806213
    lut[92] = 12'd52; // x=1.4413, y=0.808649
    lut[93] = 12'd52; // x=1.4569, y=0.811061
    lut[94] = 12'd52; // x=1.4726, y=0.813450
    lut[95] = 12'd52; // x=1.4883, y=0.815816
    lut[96] = 12'd52; // x=1.5039, y=0.818158
    lut[97] = 12'd53; // x=1.5196, y=0.820477
    lut[98] = 12'd53; // x=1.5352, y=0.822773
    lut[99] = 12'd53; // x=1.5509, y=0.825046
    lut[100] = 12'd53; // x=1.5666, y=0.827295
    lut[101] = 12'd53; // x=1.5822, y=0.829522
    lut[102] = 12'd53; // x=1.5979, y=0.831726
    lut[103] = 12'd53; // x=1.6136, y=0.833907
    lut[104] = 12'd54; // x=1.6292, y=0.836066
    lut[105] = 12'd54; // x=1.6449, y=0.838202
    lut[106] = 12'd54; // x=1.6606, y=0.840315
    lut[107] = 12'd54; // x=1.6762, y=0.842406
    lut[108] = 12'd54; // x=1.6919, y=0.844475
    lut[109] = 12'd54; // x=1.7076, y=0.846521
    lut[110] = 12'd54; // x=1.7232, y=0.848545
    lut[111] = 12'd54; // x=1.7389, y=0.850548
    lut[112] = 12'd55; // x=1.7546, y=0.852528
    lut[113] = 12'd55; // x=1.7702, y=0.854487
    lut[114] = 12'd55; // x=1.7859, y=0.856424
    lut[115] = 12'd55; // x=1.8016, y=0.858340
    lut[116] = 12'd55; // x=1.8172, y=0.860234
    lut[117] = 12'd55; // x=1.8329, y=0.862107
    lut[118] = 12'd55; // x=1.8486, y=0.863958
    lut[119] = 12'd55; // x=1.8642, y=0.865789
    lut[120] = 12'd56; // x=1.8799, y=0.867599
    lut[121] = 12'd56; // x=1.8956, y=0.869388
    lut[122] = 12'd56; // x=1.9112, y=0.871157
    lut[123] = 12'd56; // x=1.9269, y=0.872905
    lut[124] = 12'd56; // x=1.9426, y=0.874633
    lut[125] = 12'd56; // x=1.9582, y=0.876341
    lut[126] = 12'd56; // x=1.9739, y=0.878028
    lut[127] = 12'd56; // x=1.9896, y=0.879696
    lut[128] = 12'd56; // x=2.0052, y=0.881344
    lut[129] = 12'd57; // x=2.0209, y=0.882973
    lut[130] = 12'd57; // x=2.0366, y=0.884582
    lut[131] = 12'd57; // x=2.0522, y=0.886172
    lut[132] = 12'd57; // x=2.0679, y=0.887742
    lut[133] = 12'd57; // x=2.0836, y=0.889294
    lut[134] = 12'd57; // x=2.0992, y=0.890827
    lut[135] = 12'd57; // x=2.1149, y=0.892341
    lut[136] = 12'd57; // x=2.1305, y=0.893837
    lut[137] = 12'd57; // x=2.1462, y=0.895314
    lut[138] = 12'd57; // x=2.1619, y=0.896774
    lut[139] = 12'd57; // x=2.1775, y=0.898215
    lut[140] = 12'd58; // x=2.1932, y=0.899638
    lut[141] = 12'd58; // x=2.2089, y=0.901044
    lut[142] = 12'd58; // x=2.2245, y=0.902432
    lut[143] = 12'd58; // x=2.2402, y=0.903803
    lut[144] = 12'd58; // x=2.2559, y=0.905156
    lut[145] = 12'd58; // x=2.2715, y=0.906492
    lut[146] = 12'd58; // x=2.2872, y=0.907812
    lut[147] = 12'd58; // x=2.3029, y=0.909115
    lut[148] = 12'd58; // x=2.3185, y=0.910401
    lut[149] = 12'd58; // x=2.3342, y=0.911670
    lut[150] = 12'd58; // x=2.3499, y=0.912924
    lut[151] = 12'd59; // x=2.3655, y=0.914161
    lut[152] = 12'd59; // x=2.3812, y=0.915383
    lut[153] = 12'd59; // x=2.3969, y=0.916588
    lut[154] = 12'd59; // x=2.4125, y=0.917778
    lut[155] = 12'd59; // x=2.4282, y=0.918952
    lut[156] = 12'd59; // x=2.4439, y=0.920112
    lut[157] = 12'd59; // x=2.4595, y=0.921256
    lut[158] = 12'd59; // x=2.4752, y=0.922385
    lut[159] = 12'd59; // x=2.4909, y=0.923499
    lut[160] = 12'd59; // x=2.5065, y=0.924598
    lut[161] = 12'd59; // x=2.5222, y=0.925683
    lut[162] = 12'd59; // x=2.5379, y=0.926754
    lut[163] = 12'd59; // x=2.5535, y=0.927810
    lut[164] = 12'd59; // x=2.5692, y=0.928852
    lut[165] = 12'd60; // x=2.5849, y=0.929881
    lut[166] = 12'd60; // x=2.6005, y=0.930895
    lut[167] = 12'd60; // x=2.6162, y=0.931896
    lut[168] = 12'd60; // x=2.6319, y=0.932884
    lut[169] = 12'd60; // x=2.6475, y=0.933858
    lut[170] = 12'd60; // x=2.6632, y=0.934819
    lut[171] = 12'd60; // x=2.6789, y=0.935767
    lut[172] = 12'd60; // x=2.6945, y=0.936702
    lut[173] = 12'd60; // x=2.7102, y=0.937625
    lut[174] = 12'd60; // x=2.7258, y=0.938535
    lut[175] = 12'd60; // x=2.7415, y=0.939432
    lut[176] = 12'd60; // x=2.7572, y=0.940318
    lut[177] = 12'd60; // x=2.7728, y=0.941191
    lut[178] = 12'd60; // x=2.7885, y=0.942052
    lut[179] = 12'd60; // x=2.8042, y=0.942901
    lut[180] = 12'd60; // x=2.8198, y=0.943739
    lut[181] = 12'd60; // x=2.8355, y=0.944565
    lut[182] = 12'd61; // x=2.8512, y=0.945379
    lut[183] = 12'd61; // x=2.8668, y=0.946183
    lut[184] = 12'd61; // x=2.8825, y=0.946975
    lut[185] = 12'd61; // x=2.8982, y=0.947756
    lut[186] = 12'd61; // x=2.9138, y=0.948526
    lut[187] = 12'd61; // x=2.9295, y=0.949286
    lut[188] = 12'd61; // x=2.9452, y=0.950035
    lut[189] = 12'd61; // x=2.9608, y=0.950773
    lut[190] = 12'd61; // x=2.9765, y=0.951501
    lut[191] = 12'd61; // x=2.9922, y=0.952219
    lut[192] = 12'd61; // x=3.0078, y=0.952927
    lut[193] = 12'd61; // x=3.0235, y=0.953625
    lut[194] = 12'd61; // x=3.0392, y=0.954312
    lut[195] = 12'd61; // x=3.0548, y=0.954991
    lut[196] = 12'd61; // x=3.0705, y=0.955659
    lut[197] = 12'd61; // x=3.0862, y=0.956318
    lut[198] = 12'd61; // x=3.1018, y=0.956968
    lut[199] = 12'd61; // x=3.1175, y=0.957609
    lut[200] = 12'd61; // x=3.1332, y=0.958240
    lut[201] = 12'd61; // x=3.1488, y=0.958862
    lut[202] = 12'd61; // x=3.1645, y=0.959476
    lut[203] = 12'd61; // x=3.1802, y=0.960081
    lut[204] = 12'd61; // x=3.1958, y=0.960677
    lut[205] = 12'd62; // x=3.2115, y=0.961264
    lut[206] = 12'd62; // x=3.2272, y=0.961843
    lut[207] = 12'd62; // x=3.2428, y=0.962414
    lut[208] = 12'd62; // x=3.2585, y=0.962977
    lut[209] = 12'd62; // x=3.2742, y=0.963531
    lut[210] = 12'd62; // x=3.2898, y=0.964078
    lut[211] = 12'd62; // x=3.3055, y=0.964616
    lut[212] = 12'd62; // x=3.3211, y=0.965147
    lut[213] = 12'd62; // x=3.3368, y=0.965670
    lut[214] = 12'd62; // x=3.3525, y=0.966186
    lut[215] = 12'd62; // x=3.3681, y=0.966694
    lut[216] = 12'd62; // x=3.3838, y=0.967195
    lut[217] = 12'd62; // x=3.3995, y=0.967688
    lut[218] = 12'd62; // x=3.4151, y=0.968174
    lut[219] = 12'd62; // x=3.4308, y=0.968654
    lut[220] = 12'd62; // x=3.4465, y=0.969126
    lut[221] = 12'd62; // x=3.4621, y=0.969591
    lut[222] = 12'd62; // x=3.4778, y=0.970050
    lut[223] = 12'd62; // x=3.4935, y=0.970501
    lut[224] = 12'd62; // x=3.5091, y=0.970947
    lut[225] = 12'd62; // x=3.5248, y=0.971385
    lut[226] = 12'd62; // x=3.5405, y=0.971818
    lut[227] = 12'd62; // x=3.5561, y=0.972243
    lut[228] = 12'd62; // x=3.5718, y=0.972663
    lut[229] = 12'd62; // x=3.5875, y=0.973077
    lut[230] = 12'd62; // x=3.6031, y=0.973484
    lut[231] = 12'd62; // x=3.6188, y=0.973885
    lut[232] = 12'd62; // x=3.6345, y=0.974281
    lut[233] = 12'd62; // x=3.6501, y=0.974671
    lut[234] = 12'd62; // x=3.6658, y=0.975054
    lut[235] = 12'd62; // x=3.6815, y=0.975433
    lut[236] = 12'd62; // x=3.6971, y=0.975805
    lut[237] = 12'd62; // x=3.7128, y=0.976172
    lut[238] = 12'd62; // x=3.7285, y=0.976534
    lut[239] = 12'd63; // x=3.7441, y=0.976890
    lut[240] = 12'd63; // x=3.7598, y=0.977241
    lut[241] = 12'd63; // x=3.7755, y=0.977587
    lut[242] = 12'd63; // x=3.7911, y=0.977928
    lut[243] = 12'd63; // x=3.8068, y=0.978264
    lut[244] = 12'd63; // x=3.8225, y=0.978594
    lut[245] = 12'd63; // x=3.8381, y=0.978920
    lut[246] = 12'd63; // x=3.8538, y=0.979241
    lut[247] = 12'd63; // x=3.8695, y=0.979557
    lut[248] = 12'd63; // x=3.8851, y=0.979868
    lut[249] = 12'd63; // x=3.9008, y=0.980175
    lut[250] = 12'd63; // x=3.9164, y=0.980477
    lut[251] = 12'd63; // x=3.9321, y=0.980775
    lut[252] = 12'd63; // x=3.9478, y=0.981068
    lut[253] = 12'd63; // x=3.9634, y=0.981357
    lut[254] = 12'd63; // x=3.9791, y=0.981641
    lut[255] = 12'd63; // x=3.9948, y=0.981921
    lut[256] = 12'd63; // x=4.0104, y=0.982197
    lut[257] = 12'd63; // x=4.0261, y=0.982469
    lut[258] = 12'd63; // x=4.0418, y=0.982737
    lut[259] = 12'd63; // x=4.0574, y=0.983001
    lut[260] = 12'd63; // x=4.0731, y=0.983261
    lut[261] = 12'd63; // x=4.0888, y=0.983516
    lut[262] = 12'd63; // x=4.1044, y=0.983769
    lut[263] = 12'd63; // x=4.1201, y=0.984017
    lut[264] = 12'd63; // x=4.1358, y=0.984261
    lut[265] = 12'd63; // x=4.1514, y=0.984502
    lut[266] = 12'd63; // x=4.1671, y=0.984739
    lut[267] = 12'd63; // x=4.1828, y=0.984973
    lut[268] = 12'd63; // x=4.1984, y=0.985203
    lut[269] = 12'd63; // x=4.2141, y=0.985430
    lut[270] = 12'd63; // x=4.2298, y=0.985653
    lut[271] = 12'd63; // x=4.2454, y=0.985873
    lut[272] = 12'd63; // x=4.2611, y=0.986089
    lut[273] = 12'd63; // x=4.2768, y=0.986303
    lut[274] = 12'd63; // x=4.2924, y=0.986513
    lut[275] = 12'd63; // x=4.3081, y=0.986720
    lut[276] = 12'd63; // x=4.3238, y=0.986923
    lut[277] = 12'd63; // x=4.3394, y=0.987124
    lut[278] = 12'd63; // x=4.3551, y=0.987322
    lut[279] = 12'd63; // x=4.3708, y=0.987516
    lut[280] = 12'd63; // x=4.3864, y=0.987708
    lut[281] = 12'd63; // x=4.4021, y=0.987897
    lut[282] = 12'd63; // x=4.4178, y=0.988082
    lut[283] = 12'd63; // x=4.4334, y=0.988266
    lut[284] = 12'd63; // x=4.4491, y=0.988446
    lut[285] = 12'd63; // x=4.4648, y=0.988623
    lut[286] = 12'd63; // x=4.4804, y=0.988798
    lut[287] = 12'd63; // x=4.4961, y=0.988970
    lut[288] = 12'd63; // x=4.5117, y=0.989140
    lut[289] = 12'd63; // x=4.5274, y=0.989307
    lut[290] = 12'd63; // x=4.5431, y=0.989471
    lut[291] = 12'd63; // x=4.5587, y=0.989633
    lut[292] = 12'd63; // x=4.5744, y=0.989793
    lut[293] = 12'd63; // x=4.5901, y=0.989950
    lut[294] = 12'd63; // x=4.6057, y=0.990105
    lut[295] = 12'd63; // x=4.6214, y=0.990257
    lut[296] = 12'd63; // x=4.6371, y=0.990407
    lut[297] = 12'd63; // x=4.6527, y=0.990555
    lut[298] = 12'd63; // x=4.6684, y=0.990700
    lut[299] = 12'd63; // x=4.6841, y=0.990843
    lut[300] = 12'd63; // x=4.6997, y=0.990984
    lut[301] = 12'd63; // x=4.7154, y=0.991123
    lut[302] = 12'd63; // x=4.7311, y=0.991260
    lut[303] = 12'd63; // x=4.7467, y=0.991395
    lut[304] = 12'd63; // x=4.7624, y=0.991527
    lut[305] = 12'd63; // x=4.7781, y=0.991658
    lut[306] = 12'd63; // x=4.7937, y=0.991787
    lut[307] = 12'd63; // x=4.8094, y=0.991913
    lut[308] = 12'd63; // x=4.8251, y=0.992038
    lut[309] = 12'd63; // x=4.8407, y=0.992161
    lut[310] = 12'd64; // x=4.8564, y=0.992282
    lut[311] = 12'd64; // x=4.8721, y=0.992401
    lut[312] = 12'd64; // x=4.8877, y=0.992518
    lut[313] = 12'd64; // x=4.9034, y=0.992633
    lut[314] = 12'd64; // x=4.9191, y=0.992747
    lut[315] = 12'd64; // x=4.9347, y=0.992859
    lut[316] = 12'd64; // x=4.9504, y=0.992969
    lut[317] = 12'd64; // x=4.9661, y=0.993078
    lut[318] = 12'd64; // x=4.9817, y=0.993185
    lut[319] = 12'd64; // x=4.9974, y=0.993290
    lut[320] = 12'd64; // x=5.0131, y=0.993393
    lut[321] = 12'd64; // x=5.0287, y=0.993495
    lut[322] = 12'd64; // x=5.0444, y=0.993596
    lut[323] = 12'd64; // x=5.0601, y=0.993695
    lut[324] = 12'd64; // x=5.0757, y=0.993792
    lut[325] = 12'd64; // x=5.0914, y=0.993888
    lut[326] = 12'd64; // x=5.1070, y=0.993983
    lut[327] = 12'd64; // x=5.1227, y=0.994075
    lut[328] = 12'd64; // x=5.1384, y=0.994167
    lut[329] = 12'd64; // x=5.1540, y=0.994257
    lut[330] = 12'd64; // x=5.1697, y=0.994346
    lut[331] = 12'd64; // x=5.1854, y=0.994433
    lut[332] = 12'd64; // x=5.2010, y=0.994519
    lut[333] = 12'd64; // x=5.2167, y=0.994604
    lut[334] = 12'd64; // x=5.2324, y=0.994688
    lut[335] = 12'd64; // x=5.2480, y=0.994770
    lut[336] = 12'd64; // x=5.2637, y=0.994851
    lut[337] = 12'd64; // x=5.2794, y=0.994930
    lut[338] = 12'd64; // x=5.2950, y=0.995009
    lut[339] = 12'd64; // x=5.3107, y=0.995086
    lut[340] = 12'd64; // x=5.3264, y=0.995162
    lut[341] = 12'd64; // x=5.3420, y=0.995237
    lut[342] = 12'd64; // x=5.3577, y=0.995310
    lut[343] = 12'd64; // x=5.3734, y=0.995383
    lut[344] = 12'd64; // x=5.3890, y=0.995454
    lut[345] = 12'd64; // x=5.4047, y=0.995525
    lut[346] = 12'd64; // x=5.4204, y=0.995594
    lut[347] = 12'd64; // x=5.4360, y=0.995662
    lut[348] = 12'd64; // x=5.4517, y=0.995729
    lut[349] = 12'd64; // x=5.4674, y=0.995795
    lut[350] = 12'd64; // x=5.4830, y=0.995860
    lut[351] = 12'd64; // x=5.4987, y=0.995925
    lut[352] = 12'd64; // x=5.5144, y=0.995988
    lut[353] = 12'd64; // x=5.5300, y=0.996050
    lut[354] = 12'd64; // x=5.5457, y=0.996111
    lut[355] = 12'd64; // x=5.5614, y=0.996171
    lut[356] = 12'd64; // x=5.5770, y=0.996230
    lut[357] = 12'd64; // x=5.5927, y=0.996289
    lut[358] = 12'd64; // x=5.6084, y=0.996346
    lut[359] = 12'd64; // x=5.6240, y=0.996403
    lut[360] = 12'd64; // x=5.6397, y=0.996459
    lut[361] = 12'd64; // x=5.6554, y=0.996513
    lut[362] = 12'd64; // x=5.6710, y=0.996567
    lut[363] = 12'd64; // x=5.6867, y=0.996621
    lut[364] = 12'd64; // x=5.7023, y=0.996673
    lut[365] = 12'd64; // x=5.7180, y=0.996725
    lut[366] = 12'd64; // x=5.7337, y=0.996775
    lut[367] = 12'd64; // x=5.7493, y=0.996825
    lut[368] = 12'd64; // x=5.7650, y=0.996874
    lut[369] = 12'd64; // x=5.7807, y=0.996923
    lut[370] = 12'd64; // x=5.7963, y=0.996971
    lut[371] = 12'd64; // x=5.8120, y=0.997018
    lut[372] = 12'd64; // x=5.8277, y=0.997064
    lut[373] = 12'd64; // x=5.8433, y=0.997109
    lut[374] = 12'd64; // x=5.8590, y=0.997154
    lut[375] = 12'd64; // x=5.8747, y=0.997198
    lut[376] = 12'd64; // x=5.8903, y=0.997242
    lut[377] = 12'd64; // x=5.9060, y=0.997284
    lut[378] = 12'd64; // x=5.9217, y=0.997326
    lut[379] = 12'd64; // x=5.9373, y=0.997368
    lut[380] = 12'd64; // x=5.9530, y=0.997409
    lut[381] = 12'd64; // x=5.9687, y=0.997449
    lut[382] = 12'd64; // x=5.9843, y=0.997488
    lut[383] = 12'd64; // x=6.0000, y=0.997527
end

assign out = lut[in];
endmodule
